package shared_pkg;

int error_count,correct_count;
bit test_finished;

endpackage